module CPU_Controltb;
  reg[31:0] Instruct;
  reg PC,IRQ;
  wire[25:0] JT;
  wire[15:0] Imm16;
  wire[4:0] Shamt, Rd, Rt, Rs;
  wire[2:0] PCSrc;
  wire[1:0] RegDst, MemToReg;
  wire[5:0] ALUFun;
  wire RegWr,ALUSrc1,ALUSrc2,Sign,MemWr,MemRd,EXTOp,LUOp;
  CPU_Control Con(Instruct,PC,IRQ,JT,Imm16,Shamt,Rd,Rt,Rs,
                   PCSrc,RegDst,RegWr,ALUSrc1,ALUSrc2,ALUFun,
                   Sign,MemWr,MemRd,MemToReg,EXTOp,LUOp);
  initial begin
    PC=1'b0;
    IRQ=1'b0;
    Instruct=32'b000000_01111_00011_10010_00000_100000; //and
    #100 Instruct=32'b000000_01111_00011_10010_00000_100001; //andu
    #100 Instruct=32'b000000_01111_00011_10010_00000_100010; //sub
    #100 Instruct=32'b000000_01111_00011_10010_00000_100011; //subu
    #100 Instruct=32'b000000_01111_00011_10010_00000_100100; //and
    #100 Instruct=32'b000000_01111_00011_10010_00000_100101; //or
    #100 Instruct=32'b000000_01111_00011_10010_00000_100110; //xor
    #100 Instruct=32'b000000_01111_00001_10000_00000_100111; //nor
    #100 Instruct=32'b000000_00000_00011_10010_00001_000000; //sll
    #100 Instruct=32'b000000_00000_00011_10010_00001_000010; //srl
    #100 Instruct=32'b000000_00000_00011_10010_00001_000011; //sra
    #100 Instruct=32'b000000_01111_00011_10010_00000_101010; //slt
    #100 Instruct=32'b000000_01111_00000_00000_00100_001000; //jr
    #100 Instruct=32'b000000_01111_00000_01100_00100_001001; //jalr
    #100 Instruct=32'b001000_01111_00011_10010_00110_100010; //addi
    #100 Instruct=32'b001001_01111_00011_10010_11000_100010; //addiu
    #100 Instruct=32'b001100_01111_00011_10010_10101_110110; //andi
    #100 Instruct=32'b001010_01111_00011_10010_00000_100010; //slti
    #100 Instruct=32'b001011_01111_00011_10010_00000_100010; //sltiu
    #100 Instruct=32'b100011_01111_00000_00000_00100_001000; //lw
    #100 Instruct=32'b101011_01111_00000_00000_00100_001000; //sw
    #100 Instruct=32'b001111_00000_01100_01100_00100_001000; //lui
    #100 Instruct=32'b000100_01111_00011_10010_00000_100010; //beq
    #100 Instruct=32'b000101_01111_00011_10010_00000_100010; //bne
    #100 Instruct=32'b000110_01111_00000_10010_00000_100010; //blez
    #100 Instruct=32'b000111_01111_00000_10010_00000_100010; //bgtz
    #100 Instruct=32'b000001_01111_00000_10010_00000_100010; //bltz
    #100 Instruct=32'b000010_01111_00011_10010_00000_100010; //j
    #100 Instruct=32'b000011_01111_00011_10010_00000_100010; //jal
    #100 Instruct=32'b000000_00000_00000_00000_00000_000000; //nop
    #100 Instruct=32'b111111_11111_11111_11111_11111_111111; //error_instruct
    #100 IRQ=1'b1;
    #100 PC=1'b1;
  end
endmodule