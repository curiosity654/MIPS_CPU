module CPU_Instruction_Memorg(reset,PC,Instruct);
input[7:0] PC;  //only require PC[31] & PC[8:2]
input reset;
output reg[31:0] Instruct;
always@(*) 
 begin
	if(reset) Instruct<=32'b0;
	else 
	 begin
		case(PC)
		 //Software decoding:
		 8'b0_0000000: Instruct<=32'b001001_00000_01000_0000000001000000; //addiu $t0, $zero, 64
		 8'b0_0000001: Instruct<=32'b101011_00000_01000_0000000000000000; //sw    $t0, 0($zero)
		 8'b0_0000010: Instruct<=32'b001001_00000_01000_0000000001111001; //addiu $t0, $zero, 121
		 8'b0_0000011: Instruct<=32'b101011_00000_01000_0000000000000100; //sw    $t0, 4($zero)
		 8'b0_0000100: Instruct<=32'b001001_00000_01000_0000000000100100; //addiu $t0, $zero, 36
		 8'b0_0000101: Instruct<=32'b101011_00000_01000_0000000000001000; //sw    $t0, 8($zero)
		 8'b0_0000110: Instruct<=32'b001001_00000_01000_0000000000110000; //addiu $t0, $zero, 48
		 8'b0_0000111: Instruct<=32'b101011_00000_01000_0000000000001100; //sw    $t0, 12($zero)
		 8'b0_0001000: Instruct<=32'b001001_00000_01000_0000000000011001; //addiu $t0, $zero, 21
		 8'b0_0001001: Instruct<=32'b101011_00000_01000_0000000000010000; //sw    $t0, 16($zero)
		 8'b0_0001010: Instruct<=32'b001001_00000_01000_0000000000010010; //addiu $t0, $zero, 18
		 8'b0_0001011: Instruct<=32'b101011_00000_01000_0000000000010100; //sw    $t0, 20($zero)
		 8'b0_0001100: Instruct<=32'b001001_00000_01000_0000000000000010; //addiu $t0, $zero, 2
		 8'b0_0001101: Instruct<=32'b101011_00000_01000_0000000000011000; //sw    $t0, 24($zero)
		 8'b0_0001110: Instruct<=32'b001001_00000_01000_0000000001111000; //addiu $t0, $zero, 120
		 8'b0_0001111: Instruct<=32'b101011_00000_01000_0000000000011100; //sw    $t0, 28($zero)
		 8'b0_0010000: Instruct<=32'b001001_00000_01000_0000000000000000; //addiu $t0, $zero, 0
		 8'b0_0010001: Instruct<=32'b101011_00000_01000_0000000000100000; //sw    $t0, 32($zero)
		 8'b0_0010010: Instruct<=32'b001001_00000_01000_0000000000010000; //addiu $t0, $zero, 16
		 8'b0_0010011: Instruct<=32'b101011_00000_01000_0000000000100100; //sw    $t0, 36($zero)
		 8'b0_0010100: Instruct<=32'b001001_00000_01000_0000000000001000; //addiu $t0, $zero, 8
		 8'b0_0010101: Instruct<=32'b101011_00000_01000_0000000000101000; //sw    $t0, 40($zero)
		 8'b0_0010110: Instruct<=32'b001001_00000_01000_0000000000000011; //addiu $t0, $zero, 3
		 8'b0_0010111: Instruct<=32'b101011_00000_01000_0000000000101100; //sw    $t0, 44($zero)
		 8'b0_0011000: Instruct<=32'b001001_00000_01000_0000000001000110; //addiu $t0, $zero, 70
		 8'b0_0011001: Instruct<=32'b101011_00000_01000_0000000000110000; //sw    $t0, 48$(zero)
		 8'b0_0011010: Instruct<=32'b001001_00000_01000_0000000000100001; //addiu $t0, $zero, 33
		 8'b0_0011011: Instruct<=32'b101011_00000_01000_0000000000110100; //sw    $t0, 52($zero)
		 8'b0_0011100: Instruct<=32'b001001_00000_01000_0000000000000110; //addiu $t0, $zero, 6
		 8'b0_0011101: Instruct<=32'b101011_00000_01000_0000000000111000; //sw    $t0, 56($zero)
		 8'b0_0011110: Instruct<=32'b001001_00000_01000_0000000000001110; //addiu $t0, $zero, 14
		 8'b0_0011111: Instruct<=32'b101011_00000_01000_0000000000111100; //sw    $t0, 60($zero)
		 //Initial v0=1
		 8'b0_0100000: Instruct<=32'b001001_00000_00010_0000000000000001; //addiu $v0, $zero, 1       //$v0:AN
		 //record the two 4bits numbers
		 8'b0_0100001: Instruct<=32'b000000_00000_00000_0000000000000000;   //nop
		 8'b0_0100010: Instruct<=32'b100011_10000_10001_0000000000010000;   //lw   $s1, 16($s0)        //$s1:switch
		 8'b0_0100011: Instruct<=32'b000000_00000_10001_10010_00100_000010; //srl  $s2, $s1, 4	        //$s2:switch[7:4],num1
		 8'b0_0100100: Instruct<=32'b001100_10001_10001_0000000000001111;   //andi $s1, $s1, 15        //$s1:switch[3:0],num2
		 8'b0_0100101: Instruct<=32'b000000_00000_10001_01001_00000_100000; //add  $t1, $s1, $zero
		 8'b0_0100110: Instruct<=32'b000000_00000_10010_01010_00000_100000; //add  $t2, $s2, $zero
		 8'b0_0100111: Instruct<=32'b000100_01001_00000_0000000000001000;   //beq  $t1, $zero, caseC   //num1==0,result=num2
		 8'b0_0101000: Instruct<=32'b000100_01010_00000_0000000000001001;   //beq  $t2, $zero, caseD   //num2==0,result=num1
	  	//Loop1:
		 8'b0_0101001: Instruct<=32'b000100_01001_01010_0000000000001000;   //beq  $t1, $t2, caseD
		 8'b0_0101010: Instruct<=32'b000000_01001_01010_01000_00000_101010; //slt  $t0, $t1, $t2
		 8'b0_0101011: Instruct<=32'b000101_01000_00000_0000000000000010;   //bne  $t0, $zero, caseB
		 //caseA:
		 8'b0_0101100: Instruct<=32'b000000_01001_01010_01001_00000_100010; //sub  $t1, $t1, $t2       //num1>num2
		 8'b0_0101101: Instruct<=32'b000010_00000000000000000000101001;     //j    Loop1
		 //caseB:
		 8'b0_0101110: Instruct<=32'b000000_01010_01001_01010_00000_100010; //sub  $t2, $t2, $t1       //num2>num1
		 8'b0_0101111: Instruct<=32'b000010_00000000000000000000101001;     //j    Loop1
		 //caseC:
		 8'b0_0110000: Instruct<=32'b000000_01010_00000_00011_00000_100000; //add  $v1, $t2, $zero     //$v1:result
		 8'b0_0110001: Instruct<=32'b000010_00000000000000000000110011;     //j    AN                  
	  	//caseD:                  
		 8'b0_0110010: Instruct<=32'b000000_01001_00000_00011_00000_100000; //add  $v1, $t1, $zero     
		 //AN:           
		 8'b0_0110011: Instruct<=32'b000000_00000_00010_01011_00001_000010; //srl  $t3, $v0, 1         
		 8'b0_0110100: Instruct<=32'b000100_01011_00000_0000000000000101;   //beq  $t3, $zero, num1     //digital:num1
		 8'b0_0110101: Instruct<=32'b000000_00000_00010_01011_00010_000010; //srl  $t3, $v0, 2
		 8'b0_0110110: Instruct<=32'b000100_01011_00000_0000000000000101;   //beq  $t3, $zero, num2     //digital:num2
		 //out:
		 8'b0_0110111: Instruct<=32'b001001_00000_00010_0000000000000001;   //addiu $v0, $zero, 1     
		 8'b0_0111000: Instruct<=32'b000000_00000_00011_10011_00010_000000; //sll   $s3, $v1, 2         //digital:result
		 8'b0_0111001: Instruct<=32'b000010_00000000000000000000111110;     //j     Output
		 //num1:
		 8'b0_0111010: Instruct<=32'b000000_00000_10001_10011_00010_000000; //sll  $s3, $s1, 2
		 8'b0_0111011: Instruct<=32'b000010_00000000000000000000111101;     //j    shift
		 //num2:
		 8'b0_0111100: Instruct<=32'b000000_00000_10010_10011_00010_000000; //sll  $s3, $s2, 2    
		 //shift:
		 8'b0_0111101: Instruct<=32'b000000_00000_00010_00010_00001_000000; //sll  $v0, $v0, 1
		 //Output:
		 8'b0_0111110: Instruct<=32'b000010_00000000000000000000111110;     //j   Output
		 8'b0_0111111: Instruct<=32'b00000000000000000000000000000000;      //nop
		 8'b0_1000000: Instruct<=32'b11111111111111111111111111111111;      //exception
		 8'b0_1000001: Instruct<=32'b000010_00000000000000000000100001;     //j   preparation
     8'b1_0000000: Instruct<=32'b000010_00000000000000000000000100;     //j   reset
     8'b1_0000001: Instruct<=32'b000010_00000000000000000000001000;     //j   ILLOP
		 8'b1_0000010: Instruct<=32'b000000_11010_00000_00000_00000_001000; //jr  XADR
	  	//reset:
		 8'b1_0000100: Instruct<=32'b001001_00000_10100_0000000000000011;   //addiu $s4, $zero, 3  //$s4:TCON=3
		 8'b1_0000101: Instruct<=32'b001111_00000_10000_0100000000000000;   //lui   $s0, 16384
		 8'b1_0000110: Instruct<=32'b101011_10000_10100_0000000000001000;   //sw    $s4, 8($s0)
		 8'b1_0000111: Instruct<=32'b000000_00000_00000_00000_00000_001000; //jr    $zero
		 //ILLOP:
		 8'b1_0001000: Instruct<=32'b101011_10000_10100_0000000000001000;   //sw   $s4, 8($s0)
		 8'b1_0001001: Instruct<=32'b100011_10011_10101_0000000000000000;   //lw   $s5, 0($s3)     
		 8'b1_0001010: Instruct<=32'b000000_00000_00010_10110_01000_000000; //sll  $s6, $v0, 8     //$s6:{AN,digital}
		 8'b1_0001011: Instruct<=32'b000000_10101_10110_10110_00000_100000; //add  $s6, $s5, $s6
     8'b1_0001100: Instruct<=32'b100011_10000_10101_0000000000010000;   //lw   $s5, 16($s0)    //$s5:led
     8'b1_0001101: Instruct<=32'b101011_10000_10110_0000000000010100;   //sw   $s6, 20($s0)
     8'b1_0001110: Instruct<=32'b101011_10000_10101_0000000000001100;   //sw   $s5, 12($s0)
		 8'b1_0001111: Instruct<=32'b000000_11111_00000_00000_00000_001000; //jr   $Ra
		 default:	Instruct<=32'b0;
		endcase
	 end
	end
endmodule